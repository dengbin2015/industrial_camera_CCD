LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY reference_frequency IS
PORT(CLK: IN STD_LOGIC;
	 ref_clock: OUT STD_LOGIC );
END;
ARCHITECTURE reference_frequency_ARCH OF reference_frequency IS
BEGIN
PROCESS(CLK)
--VARIABLE TEMP: INTEGER RANGE 0 TO 1:=0; 
--VARIABLE TEMP: INTEGER RANGE 0 TO 3:=0; 
VARIABLE TEMP: INTEGER RANGE 0 TO 7:=0; 
--VARIABLE TEMP: INTEGER RANGE 0 TO 9:=0; 
--VARIABLE TEMP: INTEGER RANGE 0 TO 11:=0; 
--VARIABLE TEMP: INTEGER RANGE 0 TO 15:=0; 
--VARIABLE TEMP: INTEGER RANGE 0 TO 17:=0;   --no data
--VARIABLE TEMP: INTEGER RANGE 0 TO 31:=0; 
BEGIN
	IF CLK'EVENT AND CLK = '0' THEN
		TEMP := TEMP + 1;
--		IF TEMP > 0 and TEMP <= 1 THEN
--		IF TEMP > 1 and TEMP <= 3 THEN
		IF TEMP > 3 and TEMP <= 7 THEN
--      IF -TEMP > 4 and TEMP <= 9 THEN
--      IF TEMP > 5 and TEMP <= 11 THEN
--		IF TEMP > 7 and TEMP <= 15 THEN
--      IF TEMP > 8 and TEMP <= 17 THEN
--      IF TEMP > 15 and TEMP <= 31 THEN
			ref_clock <= '1';
		ELSE
			ref_clock <= '0';
		END IF;
	END IF;
END PROCESS;
END reference_frequency_ARCH;